.ckt
donington national
[3161][0][0]
[0]
[1365.706278 439.071228]
[0.000000 0.000000]
[0.000000 0.000000]
[0.000000 0.000000]
[0]
[0]
[0.000000 0.000000]
[0]
[0]
[316]
[1009.393350 370.363258]
[1019.388229 369.863392]
[1029.382750 369.353515]
[1039.376688 368.827895]
[1049.370009 368.286265]
[1059.362805 367.731541]
[1069.355282 367.169022]
[1079.347579 366.602186]
[1089.339594 366.028676]
[1099.331026 365.441723]
[1109.321633 364.836360]
[1119.311624 364.217704]
[1129.301334 363.593121]
[1139.290862 362.964719]
[1149.280237 362.333143]
[1159.269587 361.701057]
[1169.258928 361.068793]
[1179.248322 360.437618]
[1189.237952 359.811346]
[1199.227795 359.189544]
[1209.217668 358.568391]
[1219.207272 357.941584]
[1229.196505 357.307084]
[1239.185580 356.669357]
[1249.174078 356.020023]
[1259.161137 355.342820]
[1269.146021 354.626091]
[1279.127615 353.854350]
[1289.105465 353.025158]
[1299.078312 352.126450]
[1309.039357 351.085877]
[1318.916008 349.396713]
[1328.474559 346.343544]
[1337.365633 341.641117]
[1345.349981 335.477402]
[1352.305417 328.143664]
[1358.054218 319.808316]
[1362.328612 310.613560]
[1364.891971 300.787823]
[1365.706278 290.654075]
[1364.873314 280.513991]
[1362.634173 270.583932]
[1359.238517 260.987046]
[1355.173875 251.650114]
[1350.936811 242.390343]
[1346.527336 233.212489]
[1341.761296 224.216937]
[1336.565875 215.464748]
[1331.034023 206.922725]
[1325.285104 198.526720]
[1319.326448 190.280204]
[1313.101408 182.235717]
[1306.582788 174.430443]
[1299.758685 166.894894]
[1292.624089 159.657140]
[1285.197926 152.723818]
[1277.522170 146.072411]
[1269.643026 139.667657]
[1261.558004 133.530387]
[1253.241760 127.717387]
[1244.680882 122.279977]
[1235.874662 117.260343]
[1226.833702 112.689770]
[1217.592838 108.551058]
[1208.190494 104.807405]
[1198.641481 101.472256]
[1188.960417 98.562086]
[1179.181167 96.019494]
[1169.329174 93.795126]
[1159.413759 91.897054]
[1149.446492 90.321858]
[1139.436362 89.086694]
[1129.393748 88.207550]
[1119.331281 87.690463]
[1109.262069 87.560673]
[1099.203264 87.865582]
[1089.168264 88.550725]
[1079.162079 89.529706]
[1069.175311 90.671945]
[1059.179328 91.739842]
[1049.157023 92.565211]
[1039.108847 93.071281]
[1029.046546 93.310429]
[1018.978027 93.308448]
[1008.909484 93.020493]
[998.851657 92.394635]
[988.828692 91.292662]
[978.867360 89.679859]
[968.972838 87.668007]
[959.183137 85.173708]
[949.551190 82.099298]
[940.104202 78.476270]
[930.858963 74.348236]
[921.815812 69.781708]
[912.977540 64.819605]
[904.340835 59.505839]
[895.837628 53.974988]
[887.324163 48.460389]
[878.745678 43.049763]
[870.119811 37.716839]
[861.445328 32.465322]
[852.721286 27.298639]
[843.955977 22.204027]
[835.148877 17.183954]
[826.275389 12.285514]
[817.205317 7.776871]
[807.793181 4.069457]
[798.039852 1.447682]
[788.054409 0.054333]
[777.993310 0.000000]
[768.036448 1.306550]
[758.337395 3.840553]
[748.955813 7.338486]
[739.862624 11.506514]
[731.033569 16.191102]
[722.483932 21.352397]
[714.254371 26.995499]
[706.372135 33.101440]
[698.868097 39.654416]
[691.667152 46.532309]
[684.634303 53.577967]
[677.739441 60.755345]
[670.965782 68.044511]
[664.236740 75.373971]
[657.435844 82.638282]
[650.472065 89.750299]
[643.310691 96.668343]
[635.904721 103.330193]
[628.198764 109.651780]
[620.193326 115.600593]
[611.919411 121.181494]
[603.426423 126.434174]
[594.773006 131.427320]
[585.978681 136.176256]
[577.044362 140.665905]
[567.930906 144.792266]
[558.630009 148.496516]
[549.154979 151.749646]
[539.504521 154.469433]
[529.725654 156.718947]
[519.837896 158.467440]
[509.853441 159.615534]
[499.810619 160.188293]
[489.744833 160.309317]
[479.675229 160.237949]
[469.605731 160.178650]
[459.536058 160.089702]
[449.466616 159.861554]
[439.400431 159.448523]
[429.343748 158.793635]
[419.308018 157.825670]
[409.307302 156.507287]
[399.356549 154.822761]
[389.470722 152.765922]
[379.664021 150.338656]
[369.946221 147.558926]
[360.332106 144.424399]
[350.837278 140.931006]
[341.475022 137.084408]
[332.262859 132.879712]
[323.195132 128.362401]
[314.246323 123.607019]
[305.375591 118.703299]
[296.544593 113.726430]
[287.735352 108.710125]
[278.931374 103.684341]
[270.118339 98.674880]
[261.286560 93.699425]
[252.412252 88.802397]
[243.410553 84.151992]
[234.169461 80.017094]
[224.572921 76.849797]
[214.622174 75.260889]
[204.579590 75.590157]
[194.762480 77.638667]
[185.380887 81.119263]
[176.573235 85.831965]
[168.397498 91.543880]
[160.893891 98.093122]
[154.137515 105.391265]
[148.181750 113.342123]
[142.642433 121.586307]
[136.928683 129.712316]
[131.007458 137.693126]
[125.086760 145.674319]
[119.178694 153.664650]
[113.275720 161.658654]
[107.392286 169.666705]
[101.527623 177.688190]
[95.675384 185.718529]
[89.837115 193.758789]
[84.012926 201.809014]
[78.196006 209.864369]
[72.378099 217.919028]
[66.547626 225.964807]
[60.700361 233.998684]
[54.839376 242.022792]
[48.962186 250.035321]
[43.078645 258.043299]
[37.219360 266.068608]
[31.404371 274.125308]
[25.628636 282.209536]
[19.899864 290.326306]
[14.243117 298.492223]
[8.865304 306.838621]
[4.375254 315.674106]
[1.313180 325.083882]
[-0.000000 334.874631]
[0.555250 344.732927]
[2.679946 354.378453]
[6.044153 363.668022]
[10.465554 372.507653]
[15.845924 380.804404]
[22.092482 388.478867]
[29.075147 395.501583]
[36.682674 401.854404]
[44.844666 407.492370]
[53.477055 412.399368]
[62.481244 416.607963]
[71.702484 420.338992]
[81.048498 423.757056]
[90.543967 426.751982]
[100.187561 429.256100]
[109.934096 431.353260]
[119.743648 433.156460]
[129.597170 434.723294]
[139.486695 436.067380]
[149.407694 437.184382]
[159.355086 438.072302]
[169.326198 438.696078]
[179.315433 439.030181]
[189.314394 439.071228]
[199.314852 438.837099]
[209.312315 438.422353]
[219.307997 437.946104]
[229.304121 437.483742]
[239.301609 437.068462]
[249.300440 436.709213]
[259.300287 436.404979]
[269.300832 436.154299]
[279.301735 435.946049]
[289.302758 435.761453]
[299.303829 435.593064]
[309.304922 435.441229]
[319.306011 435.305636]
[329.307067 435.186583]
[339.308071 435.082532]
[349.309029 434.988393]
[359.309945 434.901775]
[369.310810 434.823168]
[379.311611 434.753331]
[389.312349 434.691298]
[399.313047 434.633946]
[409.313708 434.580625]
[419.314226 434.541383]
[429.314407 434.529914]
[439.314221 434.543509]
[449.313837 434.569161]
[459.313378 434.599084]
[469.312872 434.631721]
[479.312270 434.669578]
[489.311497 434.716544]
[499.310626 434.768525]
[509.309969 434.809269]
[519.309909 434.814184]
[529.310447 434.772571]
[539.311254 434.701826]
[549.312087 434.627755]
[559.312811 434.567214]
[569.313274 434.532847]
[579.313580 434.512038]
[589.313880 434.491704]
[599.313986 434.485793]
[609.313744 434.502791]
[619.313196 434.537689]
[629.312351 434.588275]
[639.311477 434.640350]
[649.311903 434.483748]
[659.237764 433.226940]
[668.579848 429.614750]
[676.405606 423.296589]
[682.576661 415.276286]
[688.484422 407.046758]
[695.252055 399.531382]
[702.987674 393.048467]
[711.512802 387.674680]
[720.587426 383.328860]
[730.031328 379.893872]
[739.745803 377.386563]
[749.629684 375.721529]
[759.545631 374.271592]
[769.480439 372.983365]
[779.458827 372.173835]
[789.455894 371.762561]
[799.456556 371.666931]
[809.453356 371.807927]
[819.445287 372.089444]
[829.435055 372.419392]
[839.424843 372.748945]
[849.416291 373.041914]
[859.410169 373.275313]
[869.406334 373.442561]
[879.404462 373.538947]
[889.404102 373.561940]
[899.404597 373.524139]
[909.405402 373.453667]
[919.406343 373.362128]
[929.407405 373.239284]
[939.408451 373.066783]
[949.409149 372.832428]
[959.409101 372.535386]
[969.407994 372.179065]
[979.405681 371.771203]
[989.402311 371.325264]
[999.398142 370.853638]
[1009.393350 370.363258]
