.ckt
charlotte_fullroadcourse
[3489][0][0]
[0]
[919.133310 536.665067]
[0.000000 0.000000]
[0.000000 0.000000]
[0.000000 0.000000]
[0]
[0]
[0.000000 0.000000]
[0]
[0]
[348]
[463.921211 7.281256]
[474.453523 6.158943]
[484.992614 5.094662]
[495.537641 4.083780]
[506.090003 3.143056]
[516.650524 2.286285]
[527.220114 1.533532]
[537.800291 0.921687]
[548.389578 0.459648]
[558.985701 0.146897]
[569.586780 0.000000]
[580.190181 0.050674]
[590.784338 0.520670]
[601.247652 2.186269]
[611.168549 5.837581]
[620.106581 11.422716]
[627.813919 18.534547]
[633.962066 26.936215]
[638.686197 36.150058]
[642.843917 45.607834]
[646.522959 55.232184]
[649.268270 65.112836]
[651.224519 75.140154]
[652.510739 85.238568]
[653.114391 95.364664]
[653.060921 105.472429]
[652.310358 115.513894]
[650.763778 125.417463]
[648.418230 135.117396]
[645.348347 144.568723]
[641.527273 153.694112]
[636.918932 162.394410]
[631.504456 170.558076]
[625.473270 178.232192]
[618.857241 185.353556]
[611.623925 191.789320]
[603.866991 197.523136]
[595.622602 202.465507]
[586.938912 206.509416]
[577.922648 209.674089]
[568.690505 212.067432]
[559.315096 213.745733]
[549.855845 214.771219]
[540.356220 215.162298]
[530.856915 214.913826]
[521.399063 214.018622]
[512.007314 212.584020]
[502.649531 210.935411]
[493.280125 209.355447]
[483.889992 207.905201]
[474.478182 206.604008]
[465.033375 205.572558]
[455.541613 205.168779]
[446.073422 205.988367]
[436.832017 208.313842]
[428.044626 212.092573]
[419.936449 217.261195]
[412.569292 223.525704]
[405.998731 230.689514]
[400.325617 238.654508]
[395.581845 247.270377]
[391.776834 256.402182]
[388.768264 265.877336]
[386.419882 275.576889]
[384.751839 285.454944]
[383.864877 295.476795]
[383.960481 305.589075]
[385.501532 315.654873]
[389.171702 325.256171]
[395.317863 333.638743]
[403.464380 340.260505]
[412.684542 345.410838]
[422.377923 349.657676]
[432.353827 353.222255]
[442.530314 356.189626]
[452.839111 358.676674]
[463.232894 360.790380]
[473.677558 362.643390]
[484.140018 364.395156]
[494.603235 366.142464]
[505.062130 367.915162]
[515.514561 369.725088]
[525.957965 371.585702]
[536.392185 373.496438]
[546.817403 375.454949]
[557.233999 377.458087]
[567.643323 379.498053]
[578.045442 381.573782]
[588.444859 383.662793]
[598.848637 385.730357]
[609.255940 387.780449]
[619.662413 389.834668]
[630.069059 391.888032]
[640.485578 393.891437]
[650.920587 395.797698]
[661.378994 397.572659]
[671.904537 398.874651]
[682.498423 399.285122]
[693.076310 398.700048]
[703.551784 397.191952]
[713.830122 394.746586]
[723.745599 391.182775]
[733.210752 386.615687]
[742.235852 381.285685]
[750.776886 375.262235]
[758.858366 368.677255]
[766.589620 361.714679]
[774.037332 354.473671]
[781.141851 346.924365]
[787.502312 338.801147]
[792.558199 329.899422]
[796.067040 320.374580]
[797.874655 310.486003]
[797.700902 300.548682]
[795.566532 290.946214]
[791.647712 282.029062]
[786.155517 274.079603]
[779.378064 267.283608]
[771.657236 261.648433]
[763.322810 257.021007]
[754.572537 253.276980]
[745.613733 250.078540]
[736.601513 247.038441]
[727.657709 243.798139]
[718.988481 239.865760]
[710.909882 234.793216]
[703.627777 228.569587]
[697.292661 221.326533]
[692.317384 213.016597]
[688.948354 203.842353]
[687.102265 194.159354]
[686.873312 184.220511]
[688.612460 174.328942]
[692.381199 164.893941]
[698.032151 156.325036]
[705.294465 148.931609]
[713.631451 142.655401]
[722.591477 137.224447]
[731.928336 132.414914]
[741.534425 128.124386]
[751.383418 124.379999]
[761.514756 121.422071]
[771.897092 119.414623]
[782.433666 118.365245]
[793.032342 118.326258]
[803.587345 119.336151]
[813.991866 121.378680]
[824.112607 124.509151]
[833.791578 128.779491]
[842.926978 134.074087]
[851.419855 140.301735]
[859.334873 147.215991]
[866.677245 154.696288]
[873.305889 162.773494]
[879.403332 171.230830]
[885.098888 179.940122]
[890.297772 188.926339]
[895.022567 198.144969]
[899.358908 207.531437]
[903.333754 217.056888]
[906.932792 226.710129]
[910.137306 236.480140]
[912.917091 246.356404]
[915.215083 256.329756]
[916.992131 266.381084]
[918.232212 276.483876]
[918.940789 286.609320]
[919.133310 296.729744]
[918.818232 306.819351]
[918.007724 316.853871]
[916.744053 326.816260]
[915.105609 336.702845]
[913.156588 346.515133]
[910.909471 356.246012]
[908.317232 365.869970]
[905.353311 375.363637]
[902.027692 384.714390]
[898.351607 393.910958]
[894.343956 402.946580]
[889.999635 411.802809]
[885.286542 420.442972]
[880.186172 428.832823]
[874.708454 436.953482]
[868.864510 444.786373]
[862.665224 452.312343]
[856.137788 459.527677]
[849.308397 466.430656]
[842.198646 473.017842]
[834.821196 479.276384]
[827.185304 485.188729]
[819.312544 490.754054]
[811.227344 495.979144]
[802.947539 500.863112]
[794.487417 505.400390]
[785.857860 509.577866]
[777.070697 513.383111]
[768.144590 516.820147]
[759.101386 519.907548]
[749.960487 522.664476]
[740.736581 525.101609]
[731.442288 527.226075]
[722.090922 529.055134]
[712.694675 530.609143]
[703.262345 531.896677]
[693.802762 532.934703]
[684.324225 533.751276]
[674.834307 534.395595]
[665.338609 534.928410]
[655.839804 535.387694]
[646.338908 535.788334]
[636.836387 536.134558]
[627.332131 536.405861]
[617.826492 536.586722]
[608.320301 536.665067]
[598.814614 536.635453]
[589.310513 536.502805]
[579.808959 536.269625]
[570.310362 535.950944]
[560.814367 535.570027]
[551.319561 535.163342]
[541.824468 534.762723]
[532.328589 534.379090]
[522.831987 534.011622]
[513.334404 533.667224]
[503.835170 533.364886]
[494.333906 533.121724]
[484.830902 532.939683]
[475.326842 532.802971]
[465.822214 532.695383]
[456.317246 532.607845]
[446.812104 532.531449]
[437.306858 532.462269]
[427.801530 532.399012]
[418.296180 532.337378]
[408.790826 532.276035]
[399.285472 532.214770]
[389.780153 532.150799]
[380.274840 532.086460]
[370.769384 532.033156]
[361.263679 532.001566]
[351.757696 532.002141]
[342.251510 532.040518]
[332.745264 532.109876]
[323.239046 532.206641]
[313.732932 532.331257]
[304.226925 532.474100]
[294.720945 532.620612]
[285.215004 532.772192]
[275.709263 532.945879]
[266.203787 533.143412]
[256.698203 533.331647]
[247.192099 533.448806]
[237.686542 533.417116]
[228.185311 533.178963]
[218.694143 532.705985]
[209.220997 531.967786]
[199.773713 530.956027]
[190.357831 529.685915]
[180.981499 528.149741]
[171.651380 526.350299]
[162.373138 524.295472]
[153.160486 521.957992]
[144.034925 519.292378]
[135.022281 516.255802]
[126.138318 512.848040]
[117.386612 509.100706]
[108.772151 505.034917]
[100.314791 500.637899]
[92.048317 495.875610]
[84.009592 490.719813]
[76.221144 485.173377]
[68.696320 479.254406]
[61.458451 472.967065]
[54.523664 466.325662]
[47.927942 459.324959]
[41.718537 451.954363]
[35.900303 444.246269]
[30.459631 436.243814]
[25.404270 427.969417]
[20.767287 419.429032]
[16.573469 410.636885]
[12.829874 401.618189]
[9.526864 392.404087]
[6.695446 383.008534]
[4.365960 373.448346]
[2.533622 363.753454]
[1.214765 353.947550]
[0.384114 344.061459]
[0.000000 334.123583]
[0.077730 324.153568]
[0.632823 314.172438]
[1.683089 304.204056]
[3.254816 294.275337]
[5.338596 284.412264]
[7.922214 274.639380]
[10.991965 264.979563]
[14.529996 255.453180]
[18.533235 246.084317]
[23.005450 236.900534]
[27.929299 227.921354]
[33.296921 219.170562]
[39.105205 210.675082]
[45.326945 202.447445]
[51.919446 194.485515]
[58.820929 186.765258]
[65.989197 179.270272]
[73.394677 171.989337]
[80.987289 164.887237]
[88.729522 157.935092]
[96.613364 151.130963]
[104.631237 144.472589]
[112.787117 137.970701]
[121.091232 131.644330]
[129.522840 125.475546]
[138.066320 119.450740]
[146.727931 113.584065]
[155.518062 107.897132]
[164.447082 102.414306]
[173.527317 97.166790]
[182.759000 92.170129]
[192.109351 87.382040]
[201.544662 82.750966]
[211.046188 78.247073]
[220.604132 73.855267]
[230.219383 69.581035]
[239.893273 65.431297]
[249.622874 61.404065]
[259.400639 57.486383]
[269.221414 53.669674]
[279.085135 49.956991]
[288.993687 46.356573]
[298.949020 42.877694]
[308.951102 39.525179]
[318.997885 36.298635]
[329.090682 33.207733]
[339.230321 30.261799]
[349.416576 27.468241]
[359.651306 24.843102]
[369.933699 22.395335]
[380.259521 20.121594]
[390.624169 18.015936]
[401.023348 16.072084]
[411.452407 14.280040]
[421.908060 12.634862]
[432.386537 11.126779]
[442.883873 9.742011]
[453.396894 8.468525]
[463.921211 7.281256]
