.ckt
monza_GP
[5751][0][0]
[0]
[2210.198486 1157.490845]
[0.000000 0.000000]
[0.000000 0.000000]
[0.000000 0.000000]
[0]
[0]
[0.000000 0.000000]
[0]
[0]
[574]
[1732.573975 8.689331]
[1722.510742 8.324219]
[1712.446289 7.994507]
[1702.381104 7.697021]
[1692.314941 7.433228]
[1682.248047 7.206421]
[1672.180542 7.017944]
[1662.112671 6.856201]
[1652.044556 6.705811]
[1641.976563 6.557007]
[1631.908569 6.402710]
[1621.840698 6.237671]
[1611.772949 6.061279]
[1601.705322 5.876953]
[1591.637695 5.698853]
[1581.569580 5.547729]
[1571.501221 5.429688]
[1561.432739 5.337036]
[1551.364136 5.264404]
[1541.295410 5.211792]
[1531.226685 5.178345]
[1521.157959 5.162231]
[1511.089355 5.154175]
[1501.020630 5.142334]
[1490.951904 5.123047]
[1480.883179 5.101440]
[1470.814575 5.084595]
[1460.745850 5.073486]
[1450.677124 5.060913]
[1440.608521 5.041992]
[1430.539795 5.017334]
[1420.471069 4.989990]
[1410.402344 4.961670]
[1400.333618 4.933228]
[1390.264893 4.905762]
[1380.196289 4.883301]
[1370.127563 4.868774]
[1360.058838 4.858887]
[1349.990234 4.848145]
[1339.921509 4.833862]
[1329.852783 4.812012]
[1319.784058 4.778442]
[1309.715332 4.734375]
[1299.646729 4.681152]
[1289.578003 4.620117]
[1279.509399 4.557983]
[1269.440674 4.503662]
[1259.371948 4.458618]
[1249.303223 4.419434]
[1239.234497 4.382813]
[1229.165771 4.345459]
[1219.097168 4.304688]
[1209.028442 4.257690]
[1198.959717 4.200439]
[1188.891113 4.132080]
[1178.822510 4.051880]
[1168.753906 3.955200]
[1158.685547 3.840332]
[1148.617310 3.710571]
[1138.549072 3.571045]
[1128.480957 3.427246]
[1118.412842 3.285156]
[1108.344604 3.150269]
[1098.276367 3.019165]
[1088.208130 2.889038]
[1078.139771 2.771240]
[1068.071167 2.677368]
[1058.002563 2.613525]
[1047.933838 2.576172]
[1037.865112 2.555176]
[1027.796509 2.541016]
[1017.727783 2.519775]
[1007.659058 2.471802]
[997.590576 2.377319]
[987.522400 2.236084]
[977.454529 2.070557]
[967.386780 1.899658]
[957.318970 1.728149]
[947.251160 1.560303]
[937.183167 1.404053]
[927.115051 1.258789]
[917.046875 1.122681]
[906.978577 0.991699]
[896.910339 0.860962]
[886.842102 0.727905]
[876.774048 0.580078]
[866.706055 0.421509]
[856.638184 0.257690]
[846.570313 0.095215]
[836.501831 0.000000]
[826.469910 0.707275]
[817.036194 4.001831]
[809.752808 10.779297]
[805.519653 19.800415]
[802.798157 29.421143]
[798.370605 38.332642]
[790.753113 44.735352]
[781.156555 47.526733]
[771.099609 47.628296]
[761.121887 46.296021]
[751.334290 43.917480]
[741.701721 40.959839]
[732.117920 37.845581]
[722.523560 34.764160]
[712.896118 31.788574]
[703.206665 29.024170]
[693.438538 26.554932]
[683.590881 24.429565]
[673.675049 22.653687]
[663.710571 21.178955]
[653.710815 19.973145]
[643.683594 19.030151]
[633.638306 18.311890]
[623.581848 17.784424]
[613.518188 17.436401]
[603.451050 17.224243]
[593.382813 17.091309]
[583.314331 16.994385]
[573.245728 16.908447]
[563.177124 16.835205]
[553.108398 16.796265]
[543.040039 16.837036]
[532.974121 17.032837]
[522.918335 17.496216]
[512.883118 18.275269]
[502.871826 19.309082]
[492.884460 20.546753]
[482.923431 21.975464]
[472.998657 23.630615]
[463.126434 25.567871]
[453.317230 27.796631]
[443.576782 30.303711]
[433.912842 33.086182]
[424.337982 36.156250]
[414.868011 39.531250]
[405.515137 43.213867]
[396.296570 47.216064]
[387.208344 51.502808]
[378.240356 56.032349]
[369.411987 60.824829]
[360.732483 65.878662]
[352.216187 71.199463]
[343.882355 76.798462]
[335.763580 82.700806]
[327.891235 88.924438]
[320.248962 95.425415]
[312.805634 102.151001]
[305.561584 109.087891]
[298.537018 116.244507]
[291.730652 123.606567]
[285.149811 131.168335]
[278.792786 138.917053]
[272.640686 146.827515]
[266.694397 154.891846]
[260.956909 163.104126]
[255.430847 171.458313]
[250.124786 179.952026]
[245.044724 188.580933]
[240.202728 197.343750]
[235.608673 206.237122]
[231.271011 215.256348]
[227.196976 224.395813]
[223.366440 233.638428]
[219.769806 242.972839]
[216.391022 252.386963]
[213.209885 261.868408]
[210.228912 271.413452]
[207.459427 281.020508]
[204.899521 290.684387]
[202.537445 300.397217]
[200.383759 310.157227]
[198.449493 319.961670]
[196.721451 329.803528]
[195.160248 339.672302]
[193.723602 349.559326]
[192.366684 359.457275]
[191.036285 369.358582]
[189.696213 379.258667]
[188.351837 389.158203]
[187.030487 399.060730]
[185.746704 408.968018]
[184.494904 418.879150]
[183.265182 428.792969]
[182.050735 438.708557]
[180.843155 448.625000]
[179.631470 458.540894]
[178.406204 468.455200]
[177.161865 478.367310]
[175.905304 488.277832]
[174.653366 498.189026]
[173.422852 508.102722]
[172.223526 518.020081]
[171.068344 527.942444]
[169.959991 537.869873]
[168.877289 547.800049]
[167.798706 557.730591]
[166.710342 567.660156]
[165.612259 577.588684]
[164.510986 587.516846]
[163.403885 597.444458]
[162.290527 607.371399]
[161.181519 617.298767]
[160.091339 627.228088]
[159.024643 637.159912]
[157.977753 647.093689]
[156.939606 657.028320]
[155.897675 666.962646]
[154.844528 676.895752]
[153.753754 686.825073]
[152.533569 696.739807]
[150.693100 706.557312]
[147.106140 715.865845]
[141.134888 723.869629]
[133.206116 729.977234]
[124.162117 734.332886]
[115.206848 738.853821]
[107.429848 745.159424]
[101.234612 753.013916]
[96.421791 761.785645]
[92.728752 771.076538]
[89.860512 780.654358]
[87.214180 790.295532]
[84.434624 799.899841]
[81.511024 809.462402]
[78.537987 819.010010]
[75.492142 828.535034]
[72.283264 838.007263]
[68.880707 847.413025]
[65.348434 856.771851]
[61.753517 866.107239]
[58.122738 875.428955]
[54.494488 884.751648]
[50.896969 894.086060]
[47.320072 903.428223]
[43.733555 912.766785]
[40.114197 922.092896]
[36.457935 931.404846]
[32.750992 940.697083]
[28.985559 949.966125]
[25.180958 959.219482]
[21.364979 968.468262]
[17.587561 977.732544]
[13.911729 987.036804]
[10.370581 996.392273]
[7.028722 1005.819214]
[4.030235 1015.358093]
[1.715221 1025.078247]
[0.363264 1034.972656]
[0.000000 1044.947144]
[0.742126 1054.893066]
[2.608862 1064.686890]
[5.535809 1074.212280]
[9.541818 1083.331787]
[14.592955 1091.912720]
[20.630255 1099.827393]
[27.592899 1106.938232]
[35.328686 1113.201172]
[43.667595 1118.635620]
[52.497589 1123.231689]
[61.715553 1126.992798]
[71.206146 1130.009644]
[80.863808 1132.447021]
[90.640625 1134.357178]
[100.483398 1135.905029]
[110.343361 1137.342407]
[120.212563 1138.716064]
[130.098572 1139.965210]
[140.007416 1141.022461]
[149.933014 1141.916016]
[159.862061 1142.772095]
[169.778259 1143.759766]
[179.663498 1145.012939]
[189.521591 1146.462646]
[199.379196 1147.915649]
[209.249100 1149.284302]
[219.127335 1150.593018]
[229.011185 1151.859497]
[238.899109 1153.094727]
[248.788605 1154.317383]
[258.679932 1155.525635]
[268.577881 1156.679321]
[278.509308 1157.490845]
[288.473206 1157.460083]
[298.357208 1156.188843]
[307.937897 1153.432617]
[316.930481 1149.112183]
[325.194580 1143.498413]
[332.743073 1136.941284]
[339.577606 1129.632690]
[345.789459 1121.779175]
[351.601807 1113.619873]
[357.287720 1105.370361]
[362.933167 1097.092651]
[368.434967 1088.717896]
[373.669128 1080.171509]
[378.666901 1071.482056]
[383.604431 1062.757813]
[388.599182 1054.066650]
[393.716339 1045.447998]
[398.971252 1036.913818]
[404.346680 1028.456055]
[409.795044 1020.045654]
[415.239380 1011.632629]
[420.651855 1003.198730]
[426.052368 994.757080]
[431.449371 986.313171]
[436.827026 977.856750]
[442.185211 969.387817]
[447.539734 960.916565]
[452.899109 952.448364]
[458.262329 943.982666]
[463.627167 935.518005]
[468.998169 927.057312]
[474.377991 918.602234]
[479.765686 910.152344]
[485.156921 901.704651]
[490.545258 893.255127]
[495.939148 884.809204]
[501.366425 876.385010]
[506.869598 868.010864]
[512.494263 859.718994]
[518.241943 851.513000]
[524.080627 843.372375]
[530.013184 835.300720]
[536.056885 827.313049]
[542.205505 819.406860]
[548.440979 811.569885]
[554.747620 803.790710]
[561.131775 796.075867]
[567.588440 788.422302]
[574.096802 780.813171]
[580.641174 773.235413]
[587.207336 765.676758]
[593.796692 758.138489]
[600.407959 750.619690]
[607.038757 743.118347]
[613.696594 735.641296]
[620.382507 728.189697]
[627.084534 720.752686]
[633.789673 713.318481]
[640.492676 705.882385]
[647.201416 698.451538]
[653.933472 691.042053]
[660.700684 683.665100]
[667.501099 676.319031]
[674.326904 668.996887]
[681.174805 661.695679]
[688.047302 654.417847]
[694.945190 647.164368]
[701.865906 639.932983]
[708.804626 632.719055]
[715.756226 625.517639]
[722.718628 618.326843]
[729.688232 611.143127]
[736.663391 603.964844]
[743.639954 596.787964]
[750.617249 589.611816]
[757.600098 582.441040]
[764.585510 575.272888]
[771.568970 568.102783]
[778.550232 560.930481]
[785.535522 553.762207]
[792.529419 546.602356]
[799.529785 539.449036]
[806.532715 532.298157]
[813.536865 525.148438]
[820.538269 517.996094]
[827.537170 510.841248]
[834.545288 503.695557]
[841.580017 496.576416]
[848.651306 489.493896]
[855.749817 482.439087]
[862.852478 475.388489]
[869.935181 468.317627]
[876.981201 461.209778]
[883.987244 454.062012]
[890.962769 446.884033]
[897.924622 439.692749]
[904.889038 432.503906]
[911.860962 425.322449]
[918.844849 418.152710]
[925.845703 410.999878]
[932.864746 403.864990]
[939.900879 396.747192]
[946.950317 389.642700]
[954.015808 382.554443]
[961.159058 375.545715]
[968.433044 368.674377]
[975.988831 362.120605]
[984.154114 356.363953]
[993.012573 351.760986]
[1002.423523 348.457153]
[1012.186829 346.431763]
[1022.126221 345.787354]
[1032.080811 346.254517]
[1042.015503 347.044983]
[1051.948853 347.851685]
[1061.898804 348.414246]
[1071.864624 348.319336]
[1081.791382 347.398499]
[1091.618042 345.695862]
[1101.279663 343.211060]
[1110.690308 339.889038]
[1119.797852 335.795532]
[1128.561890 331.002686]
[1136.924438 325.531067]
[1144.850830 319.437134]
[1152.609009 313.124634]
[1160.669678 307.212463]
[1169.168701 301.957886]
[1178.057861 297.404907]
[1187.268066 293.551025]
[1196.720215 290.346191]
[1206.367432 287.800659]
[1216.157349 285.888916]
[1226.041992 284.569458]
[1235.976318 283.709412]
[1245.929443 283.118286]
[1255.892334 282.745239]
[1265.859985 282.567810]
[1275.828491 282.586060]
[1285.793945 282.802795]
[1295.755493 283.147705]
[1305.715088 283.542603]
[1315.674805 283.934204]
[1325.635132 284.309937]
[1335.596069 284.671082]
[1345.557739 285.014099]
[1355.520142 285.335571]
[1365.483398 285.631958]
[1375.447632 285.899292]
[1385.412598 286.139954]
[1395.378296 286.357544]
[1405.344238 286.556152]
[1415.310791 286.732666]
[1425.277954 286.879639]
[1435.245728 286.987305]
[1445.214111 287.046997]
[1455.182739 287.058228]
[1465.151489 287.027344]
[1475.120239 286.969482]
[1485.088989 286.895935]
[1495.057617 286.812622]
[1505.026367 286.726807]
[1514.994995 286.644897]
[1524.963745 286.574524]
[1534.932495 286.519287]
[1544.901245 286.479370]
[1554.870117 286.454346]
[1564.838867 286.440063]
[1574.807617 286.429565]
[1584.776367 286.411987]
[1594.745117 286.368591]
[1604.713867 286.287476]
[1614.682251 286.171265]
[1624.650513 286.034912]
[1634.618774 285.895386]
[1644.587036 285.755493]
[1654.555298 285.615967]
[1664.523560 285.474792]
[1674.491699 285.325806]
[1684.459717 285.169067]
[1694.427612 285.002747]
[1704.395508 284.827393]
[1714.363159 284.647400]
[1724.330933 284.463867]
[1734.298584 284.277344]
[1744.266235 284.089722]
[1754.233887 283.904968]
[1764.201538 283.721069]
[1774.169189 283.534790]
[1784.136841 283.346741]
[1794.104370 283.155396]
[1804.071899 282.961304]
[1814.039429 282.765198]
[1824.006958 282.568237]
[1833.974487 282.376221]
[1843.942139 282.193726]
[1853.910034 282.020264]
[1863.877930 281.855103]
[1873.845947 281.694763]
[1883.813965 281.536377]
[1893.782104 281.380493]
[1903.750122 281.225647]
[1913.718262 281.069702]
[1923.686279 280.912048]
[1933.654175 280.750122]
[1943.622192 280.583496]
[1953.590088 280.418945]
[1963.558228 280.263123]
[1973.526367 280.118164]
[1983.494629 279.985168]
[1993.463135 279.864624]
[2003.431641 279.753174]
[2013.400146 279.640625]
[2023.368408 279.508667]
[2033.336426 279.344299]
[2043.303955 279.152710]
[2053.271240 278.942139]
[2063.238037 278.714844]
[2073.204834 278.474609]
[2083.171143 278.216309]
[2093.136475 277.921997]
[2103.100586 277.580078]
[2113.061768 277.151855]
[2123.013916 276.545654]
[2132.939697 275.591431]
[2142.777100 273.960938]
[2152.402588 271.345093]
[2161.676270 267.658203]
[2170.459717 262.908447]
[2178.629395 257.154663]
[2186.079834 250.485779]
[2192.665039 242.952881]
[2198.250732 234.642395]
[2202.772705 225.699219]
[2206.234863 216.286377]
[2208.616455 206.537720]
[2209.917969 196.579895]
[2210.198486 186.535522]
[2209.507080 176.505859]
[2207.903564 166.576416]
[2205.456299 156.816406]
[2202.220947 147.285156]
[2198.244629 138.035278]
[2193.578125 129.111084]
[2188.241455 120.568481]
[2182.285889 112.442627]
[2175.781250 104.747559]
[2168.761230 97.518433]
[2161.292725 90.751831]
[2153.434326 84.441650]
[2145.244629 78.567017]
[2136.790039 73.079834]
[2128.114502 67.949341]
[2119.239502 63.173218]
[2110.175781 58.766113]
[2100.946533 54.717651]
[2091.570801 51.022827]
[2082.069580 47.665039]
[2072.462891 44.623535]
[2062.764893 41.889771]
[2052.991211 39.442871]
[2043.160767 37.236694]
[2033.287109 35.234985]
[2023.381470 33.399780]
[2013.451782 31.701416]
[2003.502808 30.122070]
[1993.539673 28.636841]
[1983.565308 27.229736]
[1973.581543 25.893433]
[1963.588989 24.624756]
[1953.587646 23.430176]
[1943.577637 22.312256]
[1933.560181 21.265015]
[1923.536743 20.277832]
[1913.509277 19.335205]
[1903.478271 18.431152]
[1893.444214 17.563965]
[1883.406860 16.737427]
[1873.365723 15.959595]
[1863.320313 15.240112]
[1853.271118 14.580322]
[1843.219116 13.966431]
[1833.165527 13.380981]
[1823.110718 12.819092]
[1813.054565 12.282959]
[1802.997070 11.773804]
[1792.938599 11.286377]
[1782.879517 10.809937]
[1772.820068 10.343994]
[1762.759888 9.897827]
[1752.698608 9.475952]
[1742.636475 9.076294]
