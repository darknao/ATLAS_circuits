.ckt
spa combined
[6931][0][0]
[0]
[1996.194394 1532.847049]
[0.000000 0.000000]
[0.000000 0.000000]
[0.000000 0.000000]
[0]
[0]
[0.000000 0.000000]
[0]
[0]
[693]
[1646.740606 254.398695]
[1656.002438 250.053304]
[1665.260187 245.700850]
[1674.508953 241.332902]
[1683.747342 236.947132]
[1692.973644 232.540713]
[1702.189577 228.116662]
[1711.404244 223.690461]
[1720.627038 219.278068]
[1729.862616 214.887488]
[1739.108155 210.513986]
[1748.358152 206.148155]
[1757.613017 201.790719]
[1766.878117 197.450997]
[1776.157462 193.136067]
[1785.451868 188.847526]
[1794.761842 184.586460]
[1804.086868 180.352148]
[1813.424240 176.139925]
[1822.768823 171.940664]
[1832.109569 167.734500]
[1841.434525 163.500073]
[1850.742257 159.235036]
[1860.046163 154.963229]
[1869.363903 150.715951]
[1878.704176 146.508955]
[1888.068155 142.344807]
[1897.455042 138.222543]
[1906.866119 134.145034]
[1916.301249 130.112563]
[1925.756878 126.118915]
[1935.231812 122.162215]
[1944.728955 118.248505]
[1954.242606 114.367047]
[1963.746199 110.465922]
[1973.205197 106.478833]
[1982.490097 102.176523]
[1991.229054 97.033160]
[1996.194394 89.004645]
[1992.642607 80.997423]
[1984.536850 76.728919]
[1975.879522 73.539684]
[1967.185293 70.439845]
[1958.492966 67.335317]
[1949.805515 64.218803]
[1941.121996 61.092651]
[1932.423334 58.003858]
[1923.692680 54.995227]
[1914.938903 52.045782]
[1906.164652 49.149764]
[1897.366215 46.318033]
[1888.549187 43.536608]
[1879.719353 40.790351]
[1870.876483 38.080326]
[1862.018080 35.414064]
[1853.137517 32.811411]
[1844.222534 30.310458]
[1835.265714 27.938070]
[1826.270171 25.690196]
[1817.237194 23.568613]
[1808.170110 21.567576]
[1799.076535 19.664424]
[1789.959569 17.851204]
[1780.818653 16.133857]
[1771.653574 14.517535]
[1762.468047 12.990470]
[1753.264313 11.546329]
[1744.037779 10.211281]
[1734.783223 9.019351]
[1725.497102 8.003909]
[1716.180583 7.178136]
[1706.837097 6.544646]
[1697.466605 6.139099]
[1688.071699 5.993123]
[1678.658926 6.110576]
[1669.235953 6.464584]
[1659.809014 6.992465]
[1650.381177 7.616381]
[1640.953270 8.259665]
[1631.525489 8.870372]
[1622.098053 9.434998]
[1612.671014 9.964876]
[1603.244208 10.478015]
[1593.817524 10.983267]
[1584.391296 11.462252]
[1574.966178 11.888684]
[1565.542397 12.263773]
[1556.119758 12.601490]
[1546.697936 12.914887]
[1537.276175 13.226511]
[1527.853868 13.554101]
[1518.430997 13.898923]
[1509.007556 14.262252]
[1499.583160 14.659641]
[1490.157961 15.088987]
[1480.732507 15.529411]
[1471.306889 15.977384]
[1461.881274 16.425234]
[1452.456286 16.845921]
[1443.032029 17.237842]
[1433.608852 17.592899]
[1424.190636 17.818710]
[1414.789553 17.757046]
[1405.435717 17.215881]
[1396.176887 16.056299]
[1387.077429 14.185614]
[1378.155662 11.707844]
[1369.311040 9.002700]
[1360.422115 6.425299]
[1351.444073 4.121449]
[1342.375562 2.127294]
[1333.179810 0.656620]
[1323.842774 0.000000]
[1314.425822 0.287843]
[1305.023318 1.594320]
[1295.712769 3.773195]
[1286.497130 6.484302]
[1277.368442 9.574723]
[1268.358734 13.097987]
[1259.522165 17.147241]
[1250.901509 21.746113]
[1242.525500 26.874230]
[1234.297413 32.290670]
[1225.965691 37.507270]
[1217.412806 42.261925]
[1208.794893 46.870445]
[1200.102034 51.295916]
[1191.105954 54.844988]
[1181.845468 57.310582]
[1172.489323 59.168013]
[1163.106970 60.783377]
[1153.708273 62.209571]
[1144.301858 63.528512]
[1134.894146 64.827555]
[1125.487929 66.149598]
[1116.084951 67.518907]
[1106.684925 68.928975]
[1097.284856 70.338461]
[1087.883063 71.724510]
[1078.479196 73.081280]
[1069.070816 74.369027]
[1059.657231 75.567407]
[1050.241260 76.719626]
[1040.824261 77.850343]
[1031.406197 78.957695]
[1021.987661 80.054343]
[1012.569215 81.153040]
[1003.150732 82.250903]
[993.731825 83.338890]
[984.312687 84.421392]
[974.894295 85.521263]
[965.477100 86.647761]
[956.059907 87.774332]
[946.641005 88.862107]
[937.221288 89.930549]
[927.803691 91.047760]
[918.391933 92.278085]
[908.995746 93.733020]
[899.635126 95.548816]
[890.334026 97.795428]
[881.104241 100.438151]
[871.947253 103.413158]
[862.866062 106.687365]
[853.851164 110.196432]
[844.871568 113.822499]
[835.895443 117.459778]
[826.911379 121.071408]
[817.921217 124.663173]
[808.924931 128.234830]
[799.916275 131.765368]
[790.887706 135.228354]
[781.836923 138.613891]
[772.769181 141.938721]
[763.695118 145.240547]
[754.625988 148.560349]
[745.566425 151.914687]
[736.513024 155.291033]
[727.461628 158.674496]
[718.411011 162.060715]
[709.360441 165.447102]
[700.308088 168.827169]
[691.253080 172.197802]
[682.195888 175.560641]
[673.136701 178.916344]
[664.075634 182.265304]
[655.011937 185.604792]
[645.943770 188.928109]
[636.869874 192.230538]
[627.790871 195.514207]
[618.708717 198.786224]
[609.624290 202.049807]
[600.536611 205.301258]
[591.444718 208.536904]
[582.348747 211.757160]
[573.249336 214.964355]
[564.145972 218.156442]
[555.036676 221.325685]
[545.920570 224.468429]
[536.798267 227.586800]
[527.671370 230.686934]
[518.543486 233.783134]
[509.419135 236.893388]
[500.299934 240.023995]
[491.184744 243.170329]
[482.071310 246.323516]
[472.957126 249.473783]
[463.840778 252.615588]
[454.721726 255.746788]
[445.599544 258.865641]
[436.473780 261.970285]
[427.343390 265.056446]
[418.206792 268.117569]
[409.063485 271.151317]
[399.914661 274.162315]
[390.762350 277.158809]
[381.608940 280.150712]
[372.456161 283.145255]
[363.304236 286.143359]
[354.153072 289.144636]
[345.002253 292.147350]
[335.849792 295.143217]
[326.692671 298.119531]
[317.527585 301.062007]
[308.352931 303.963152]
[299.169691 306.826523]
[289.980757 309.664470]
[280.787397 312.482418]
[271.586060 315.263795]
[262.374847 317.999018]
[253.158007 320.707492]
[243.939813 323.409460]
[234.719039 326.098975]
[225.492027 328.758040]
[216.256357 331.374025]
[207.008632 333.928283]
[197.744098 336.392807]
[188.481453 338.867525]
[179.320320 341.814066]
[170.700929 346.351404]
[163.178379 352.862752]
[156.995086 360.882488]
[152.805111 370.309571]
[150.642045 380.592819]
[149.992470 391.185094]
[150.044337 401.849622]
[149.134121 412.402091]
[146.310083 422.461422]
[141.683603 431.659180]
[135.549858 439.726839]
[128.019957 446.218905]
[119.539873 451.115096]
[110.692633 455.136115]
[101.730163 458.816137]
[92.705383 462.291708]
[83.646488 465.648393]
[74.574884 468.959190]
[65.498486 472.252453]
[56.426954 475.563504]
[47.382967 478.972684]
[38.476966 482.819274]
[29.958828 487.635443]
[22.164217 493.759339]
[15.462442 501.269538]
[10.313791 510.117559]
[6.878449 519.939471]
[4.774968 530.244617]
[3.755262 540.788569]
[3.725499 551.445146]
[4.300963 562.123666]
[4.991457 572.802064]
[5.521836 583.480635]
[5.851772 594.156143]
[6.035234 604.826864]
[6.101472 615.492166]
[6.076641 626.152335]
[6.001683 636.809321]
[5.898171 647.464373]
[5.776057 658.118123]
[5.641921 668.771011]
[5.491909 679.422737]
[5.321755 690.072955]
[5.137066 700.722060]
[4.954701 711.371344]
[4.779461 722.021176]
[4.589358 732.669856]
[4.362173 743.315575]
[4.094027 753.957865]
[3.786773 764.596723]
[3.440597 775.232011]
[3.057218 785.863745]
[2.639176 796.492040]
[2.181982 807.116303]
[1.654168 817.732870]
[1.013621 828.336122]
[0.334948 838.934646]
[0.000000 849.569280]
[0.827913 860.233477]
[3.851560 870.578999]
[9.378105 879.921985]
[16.684709 887.996521]
[25.301529 894.613854]
[35.126723 899.064906]
[45.620736 901.040171]
[56.167389 900.812104]
[66.215609 898.277785]
[75.242930 893.581282]
[82.926146 887.203493]
[88.509214 879.231100]
[91.617453 870.223108]
[92.812187 860.899141]
[92.590915 851.585412]
[91.420715 842.389905]
[89.738485 833.298255]
[87.825505 824.262641]
[85.927042 815.223325]
[84.166121 806.149824]
[82.502484 797.053274]
[80.834362 787.957765]
[79.155672 778.864697]
[77.508016 769.764469]
[75.824066 760.672665]
[74.117700 751.586078]
[72.744219 742.428734]
[72.379739 733.129584]
[73.658331 723.815164]
[76.949701 714.855335]
[82.129584 706.632907]
[89.028552 699.546470]
[97.361728 693.879017]
[106.522736 689.372682]
[116.085627 685.592196]
[125.786776 682.099552]
[135.479287 678.588100]
[145.111789 674.948295]
[154.687543 671.191016]
[164.228061 667.362750]
[173.749979 663.497569]
[183.266921 659.622577]
[192.779937 655.739874]
[202.278061 651.828068]
[211.752754 647.870915]
[221.209673 643.879714]
[230.652184 639.861168]
[240.065896 635.788603]
[249.439372 631.641805]
[258.768486 627.414870]
[268.036886 623.081052]
[277.229016 618.617035]
[286.350167 614.035661]
[295.423901 609.377819]
[304.471191 604.678021]
[313.500944 599.950652]
[322.526549 595.216788]
[331.560332 590.495733]
[340.597659 585.780240]
[349.625908 581.050516]
[358.638262 576.295999]
[367.633415 571.514826]
[376.609059 566.703649]
[385.561460 561.857025]
[394.489633 556.973794]
[403.393681 552.054456]
[412.277073 547.104461]
[421.155974 542.147829]
[430.047628 537.210065]
[438.953421 532.293314]
[447.870185 527.392955]
[456.801934 522.515100]
[465.749032 517.660423]
[474.700795 512.812816]
[483.652735 507.965478]
[492.614230 503.132677]
[501.613336 498.357695]
[510.742566 493.790537]
[520.154556 489.719794]
[529.982468 486.532501]
[540.195358 484.443543]
[550.651395 483.418396]
[561.231464 483.470729]
[571.818843 484.619707]
[582.298574 486.825606]
[592.557760 490.075185]
[602.493602 494.322986]
[612.039667 499.458351]
[621.142358 505.389345]
[629.769160 512.022648]
[637.906930 519.263771]
[645.647138 526.937582]
[653.194812 534.803429]
[660.682418 542.726932]
[668.166196 550.654074]
[675.594193 558.633592]
[682.741781 566.863863]
[689.354374 575.525044]
[695.239993 584.683750]
[700.287918 594.310712]
[704.575132 604.279240]
[708.250741 614.468907]
[711.362584 624.823187]
[713.876868 635.313440]
[715.717112 645.911591]
[716.802326 656.575606]
[717.080079 667.246911]
[716.586450 677.865118]
[715.400951 688.383863]
[713.571481 698.764942]
[711.165472 708.984573]
[708.232031 719.022688]
[704.778419 728.848540]
[700.864826 738.457932]
[696.622022 747.894492]
[692.156498 757.204866]
[687.535548 766.422648]
[682.815019 775.579056]
[678.041836 784.702362]
[673.260030 793.820202]
[668.495216 802.948807]
[663.750573 812.090134]
[659.024225 821.242941]
[654.316261 830.407228]
[649.630067 839.585036]
[644.968318 848.777939]
[640.317327 857.977456]
[635.650956 867.167510]
[630.953731 876.338473]
[626.226419 885.490673]
[621.472517 894.626167]
[616.690201 903.743678]
[611.870968 912.837618]
[607.008726 921.903819]
[602.107094 930.944345]
[597.175654 939.965267]
[592.219918 948.970093]
[587.244675 957.961925]
[582.258885 966.946703]
[577.267500 975.927732]
[572.272384 984.906257]
[567.274261 993.882762]
[562.283087 1002.863931]
[557.337342 1011.875353]
[552.646471 1021.048963]
[548.636233 1030.604896]
[545.740903 1040.650020]
[544.162683 1051.084049]
[543.964600 1061.723502]
[545.441376 1072.347536]
[548.663963 1082.662279]
[553.278856 1092.488134]
[558.971835 1101.762612]
[565.660209 1110.360501]
[573.393332 1118.029301]
[582.126530 1124.502091]
[591.718198 1129.523886]
[601.875072 1133.121246]
[612.208183 1136.097745]
[622.400099 1139.588306]
[632.179918 1144.210141]
[641.332459 1150.051148]
[649.686565 1157.026211]
[657.099159 1165.009819]
[663.485254 1173.831333]
[668.745450 1183.345232]
[672.824671 1193.389179]
[675.662757 1203.804330]
[677.169756 1214.433437]
[677.402528 1225.100058]
[676.472307 1235.657858]
[674.558353 1246.016000]
[672.029143 1256.196799]
[669.200598 1266.274796]
[666.235503 1276.302325]
[663.238342 1286.317643]
[660.221157 1296.325254]
[657.175891 1306.321987]
[654.135599 1316.320652]
[651.134459 1326.334432]
[648.177692 1336.365127]
[645.259461 1346.410315]
[642.351874 1356.459480]
[639.419962 1366.499545]
[636.469993 1376.532817]
[633.521641 1386.566700]
[630.561062 1396.595956]
[627.556942 1406.608587]
[624.482584 1416.593908]
[621.448514 1426.594855]
[618.992775 1436.795336]
[618.138578 1447.348826]
[619.726703 1457.947954]
[623.733504 1468.001669]
[629.860743 1476.979211]
[637.673187 1484.557064]
[646.689494 1490.601343]
[656.540076 1495.045827]
[666.744669 1498.505905]
[677.038925 1501.639517]
[687.369686 1504.625799]
[697.709497 1507.573907]
[708.046923 1510.532164]
[718.384726 1513.488816]
[728.723758 1516.440244]
[739.061490 1519.397211]
[749.408300 1522.315127]
[759.779089 1525.126368]
[770.184066 1527.775180]
[780.639894 1530.151219]
[791.176002 1531.955462]
[801.772866 1532.847049]
[812.341497 1532.720602]
[822.747369 1531.439301]
[832.809161 1528.874280]
[842.433296 1525.226553]
[851.586833 1520.705737]
[860.155183 1515.324663]
[868.033809 1509.126368]
[875.174655 1502.220117]
[881.544552 1494.709117]
[887.217808 1486.745614]
[892.381667 1478.499975]
[897.199671 1470.084565]
[901.787669 1461.565174]
[906.248070 1452.991137]
[910.592587 1444.369439]
[914.754898 1435.676224]
[918.689976 1426.899364]
[922.395215 1418.044108]
[925.872528 1409.117214]
[929.139253 1400.129297]
[932.211468 1391.089504]
[935.083982 1382.000762]
[937.742159 1372.864331]
[940.149843 1363.678407]
[942.290675 1354.446868]
[944.183974 1345.179586]
[945.849215 1335.884957]
[947.290281 1326.568632]
[948.512317 1317.235972]
[949.539314 1307.892797]
[950.380634 1298.543221]
[951.038318 1289.190657]
[951.550245 1279.838069]
[951.957442 1270.486804]
[952.276166 1261.137521]
[952.518620 1251.790569]
[952.687326 1242.446443]
[952.756064 1233.107041]
[952.690469 1223.775548]
[952.472474 1214.455201]
[952.100672 1205.148459]
[951.570712 1195.858232]
[950.869371 1186.588769]
[949.945649 1177.350886]
[948.728708 1168.162374]
[947.214655 1159.032845]
[945.421874 1149.967346]
[943.356709 1140.972532]
[941.029578 1132.053537]
[938.483763 1123.203643]
[935.781315 1114.406726]
[932.962420 1105.651073]
[930.078095 1096.919306]
[927.178065 1088.193351]
[924.293729 1079.461586]
[921.446936 1070.716036]
[918.647805 1061.953223]
[915.891928 1053.174975]
[913.169702 1044.384873]
[910.464007 1035.588994]
[907.761094 1026.792146]
[905.067457 1017.992078]
[902.403166 1009.181892]
[899.794377 1000.352847]
[897.265024 991.497433]
[894.868326 982.599702]
[892.684459 973.638257]
[890.743872 964.610018]
[888.985932 955.535772]
[887.337265 946.435808]
[885.815220 937.307780]
[884.525020 928.132923]
[883.596816 918.896191]
[883.112550 909.601733]
[883.081016 900.268794]
[883.494801 890.918216]
[884.329423 881.568960]
[885.529164 872.235202]
[887.079959 862.929208]
[888.990963 853.664577]
[891.256302 844.453627]
[893.866919 835.307546]
[896.812845 826.236612]
[900.093660 817.252978]
[903.695320 808.364622]
[907.571741 799.567193]
[911.638165 790.837754]
[915.823245 782.153076]
[920.094909 773.502151]
[924.394625 764.862344]
[928.643692 756.202526]
[932.812842 747.511708]
[936.931893 738.801839]
[941.035246 730.086067]
[945.129299 721.366816]
[949.210882 712.642915]
[953.298892 703.921409]
[957.427735 695.215248]
[961.668312 686.552203]
[966.134433 677.980959]
[970.907787 669.545002]
[976.068552 661.298005]
[981.792707 653.365248]
[988.189262 645.872011]
[995.195000 638.848109]
[1002.744824 632.313449]
[1010.793591 626.296946]
[1019.273659 620.795561]
[1028.136515 615.818462]
[1037.326447 611.353147]
[1046.737938 607.277356]
[1056.284624 603.461971]
[1065.935435 599.861089]
[1075.656600 596.412688]
[1085.408492 593.033122]
[1095.163881 589.661480]
[1104.909837 586.268476]
[1114.646474 582.854493]
[1124.375989 579.424566]
[1134.097451 575.976702]
[1143.807377 572.503308]
[1153.503700 569.000046]
[1163.188217 565.471065]
[1172.868123 561.932086]
[1182.553094 558.404089]
[1192.248721 554.899304]
[1201.953162 551.413826]
[1211.658108 547.929458]
[1221.356666 544.431079]
[1231.044980 540.910349]
[1240.702184 537.322731]
[1250.291270 533.592946]
[1259.791413 529.685415]
[1269.199310 525.602308]
[1278.500502 521.326212]
[1287.678625 516.839054]
[1296.726751 512.141050]
[1305.653086 507.255333]
[1314.472404 502.212031]
[1323.183524 497.015747]
[1331.784661 491.669903]
[1340.289053 486.197072]
[1348.723628 480.635129]
[1357.115694 475.019942]
[1365.492578 469.385913]
[1373.880452 463.765511]
[1382.290010 458.172121]
[1390.720614 452.605132]
[1399.174423 447.067472]
[1407.650043 441.557574]
[1416.142828 436.069671]
[1424.654363 430.605944]
[1433.193582 425.178201]
[1441.763467 419.790694]
[1450.364327 414.444277]
[1459.006294 409.153086]
[1467.707467 403.942884]
[1476.457827 398.801145]
[1484.985852 393.363038]
[1491.496241 386.064565]
[1491.291012 377.133027]
[1484.823744 370.802790]
[1477.637103 365.189485]
[1472.390892 357.755625]
[1470.494435 348.802335]
[1473.370896 339.831318]
[1480.244658 332.772473]
[1488.802513 327.375751]
[1497.839225 322.662957]
[1507.137177 318.381516]
[1516.511749 314.236658]
[1525.840780 310.009768]
[1535.091825 305.645894]
[1544.307078 301.220687]
[1553.544456 296.833256]
[1562.822021 292.515247]
[1572.133949 288.257681]
[1581.480746 284.062448]
[1590.847039 279.902491]
[1600.211913 275.739954]
[1609.559068 271.545354]
[1618.881674 267.306737]
[1628.183706 263.031633]
[1637.469690 258.728311]
[1646.740606 254.398695]
